//lesson01_top.v
//Material del Workshop: "Como crear tu propio juego Arcade (y sobrevivir al intento)"
module lesson01_top (
  input wire clk,
  input wire reset
  //output wire [3:0] video_r,
  //output wire [3:0] video_g,
  //output wire [3:0] video_b,
  //output wire csync
);
  
  //Vamos a crear un circuito con dos interruptores como entrada,
  //Vamos a aplicar varias puertas logicas a estas entradas y ver que 
  //salida producen
  
  

endmodule
  
